Name,Type,KindNO_CHIP,+def,CMD_LINE definesMOD_DIS,+def,CMD_LINE definesUSER_TEST,test,PlusargTEST,value,PlusargVSIM_TB,+def,TB definesDQ_IQP,+def,TB definesNCVERILOG,+def,TB definesjss_m10,+def,TB definestt_110,+def,TB defines