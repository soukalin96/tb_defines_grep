`ifdef VSIM_TB
`ifndef NO_CHIP
`elsif MOD_DIS