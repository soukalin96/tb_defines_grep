`ifdef VSIM_TB
`ifdef VSIM_TB
`ifdef VSIM_TB
`ifndef NO_CHIP
`elsif MOD_DIS
`ifdef DQ_IQP
`ifdef NCVERILOG

`ifdef jss_m10
`ifdef tt_110
