`define PATH top.tb.a.b.c
`define PATH2 top.tb.a.b.c
`define master(ARG) asdas
`define STACK 8
`define massster2(SID, PC, BA) asd\
`define STACKYO
