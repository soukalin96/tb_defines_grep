`define PATH top.tb.a.b.c
`define PATH2 top.tb.a.b.c
`define master(ARG) x.y.z``ARG```.a.b.c
`define STACK 8
`define master2(ARG) yolo```Mate```